`timescale 1ns / 1ps
module tb_xor_gate;
    reg a, b;
    wire y;

    xor_gate uut(a, b, y);

    initial begin
        $dumpfile("xor_gate.vcd");
        $dumpvars(0, tb_xor_gate);
        $display("A B | Y");
        $display("-------");

        a=0; b=0; #10; $display("%b %b | %b", a, b, y);
        a=0; b=1; #10; $display("%b %b | %b", a, b, y);
        a=1; b=0; #10; $display("%b %b | %b", a, b, y);
        a=1; b=1; #10; $display("%b %b | %b", a, b, y);
        $finish;
    end
endmodule
