
module not_gate(input a, output y);
    assign y = ~a;
endmodule

