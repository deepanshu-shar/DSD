`timescale 1ns / 1ps
module not_gate(input a, output y);
    assign y = ~a;
endmodule
